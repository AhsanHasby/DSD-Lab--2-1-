module RippleAdder(S, Cout, A, B, Cin);
input [3:0]A, B;
input Cin;
output [3:0]S;
output Cout;
wire [3:1]C;
FullAdder fa0(S[0], C[1], A[0], B[0], Cin);
FullAdder fa1(S[1], C[2], A[1], B[1], C[1]);
FullAdder fa2(S[2], C[3], A[2], B[2], C[2]);
FullAdder fa3(S[3], Cout, A[3], B[3], C[3]);
endmodule

module AddSub(S, Cout, A, B, mode);
input [3:0] A, B;
input mode;
output [3:0] S;
output Cout;
wire [3:0] D;
xor(D[0], B[0], mode);
xor(D[1], B[1], mode);
xor(D[2], B[2], mode);
xor(D[3], B[3], mode);
RippleAdder R1(S, Cout, A, D, mode);
endmodule


module simulate;
reg [3:0] A, B;
reg mode;
wire [3:0] S;
wire Cout;
AddSub AS1(S, Cout, A, B, mode);
initial
begin
     	A=4'b0101; B=4'b1110; mode = 1'b0;
#50	A=4'b0110; B=4'b0010; mode = 1'b0;
#50	A=4'b0101; B=4'b1110; mode = 1'b1;
#50	A=4'b0110; B=4'b0010; mode = 1'b1;

end
endmodule